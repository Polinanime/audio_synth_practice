`timescale 1ns/1ps
`define AUDIO_SQUARE
`include "../utils/test.sv"

module tb_audio_square;
  tb_audio tb();
endmodule