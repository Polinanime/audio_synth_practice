`timescale 1ns/1ps
`define AUDIO_SAW_INV
`include "../utils/test.sv"

module tb_audio_saw_inv;
  tb_audio tb();
endmodule