`timescale 1ns/1ps
`define AUDIO_NOISE
`include "../utils/test.sv"

module tb_audio_noise;
tb_audio tb();
endmodule