`timescale 1ns/1ps
`define AUDIO_SINE
`include "../utils/test.sv"

module tb_audio_sine;
tb_audio tb();
endmodule