`timescale 1ns/1ps
`define AUDIO_TRIANGLE
`include "../utils/test.sv"

module tb_audio_triangle;
tb_audio tb();
endmodule