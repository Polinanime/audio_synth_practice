`timescale 1ns/1ps
`define AUDIO_SAW
`include "../utils/test.sv"

module tb_audio_saw;
  tb_audio tb();
endmodule